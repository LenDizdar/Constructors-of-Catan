Blue
1 2 1 2 3 r 16 36 19 h 10 B 15 T 27 H
0 0 1 0 3 r 11 h 44 B 20 B
0 0 0 0 0 r h
0 0 0 0 0 r h
4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 4 11 
8
