Blue
0 0 0 0 0 r h
0 0 0 0 0 r h
0 0 0 0 0 r h
0 0 0 0 0 r h
3 11 0 10 4 9 1 3 3 4 4 10 0 5 2 11 4 5 3 3 0 9 2 12 1 8 1 6 0 6 1 4 5 7 2 2 2 8 
-1
