Yellow
0 0 0 0 2 r h 28 B 4 B
0 0 0 0 0 r h 45 B 20 B
0 0 0 0 2 r h 31 B 15 B
0 0 0 0 0 r h 8 B 35 B
0 11 3 2 4 5 1 10 4 6 4 5 3 12 3 11 1 9 5 7 1 8 2 9 2 6 0 3 0 3 2 8 0 10 2 4 1 4 
11
