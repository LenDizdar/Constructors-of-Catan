Blue
100 100 100 100 100 r 66 62 h 26 T 51 B 47 B
100 100 100 100 100 r 36 40 h 14 B 28 B 33 H
100 100 100 100 100 r 23 15 h 40 B 21 B 9 H
100 100 100 100 100 r h 44 B 31 B
2 11 4 8 5 7 2 5 1 10 1 5 2 3 0 4 4 2 0 6 0 3 3 8 3 9 2 12 0 11 1 10 1 9 4 6 3 4 
2
