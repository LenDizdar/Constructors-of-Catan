Red
0 0 0 1 0 r h 19 B 10 B
0 0 0 0 0 r h 45 B 35 B
1 0 0 0 0 r h 15 B 46 B
1 0 0 0 0 r h 22 B 20 B
1 2 2 3 4 11 3 5 2 4 0 6 2 9 0 5 1 3 4 10 1 12 5 7 0 8 3 10 4 9 0 8 3 4 2 11 1 6 
-1
