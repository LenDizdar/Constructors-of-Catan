Blue
0 1 2 0 0 r h 45 B 7 B
0 0 1 0 0 r h 18 B 51 B
0 0 0 1 0 r h 9 B 43 B
0 0 0 0 0 r h 20 B 22 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
17
